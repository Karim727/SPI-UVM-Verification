package SPI_pkg_agent;
    import uvm_pkg::*;
    import SPI_sequencer_pkg::*;
    import SPI_driver_pkg::*;
    import SPI_pkg_mon::*;
    import SPI_pkg_obj::*;
    import SPI_seq_item_pkg::*;
    `include "uvm_macros.svh"
    class SPI_agent extends uvm_agent;
        `uvm_component_utils(SPI_agent)
        SPI_sequencer sqr;
        SPI_driver drv;
        SPI_mon mon;
        SPI_config_obj SPI_cfg;
        uvm_analysis_port #(SPI_seq_item) agt_ap;
        function new(string name = "SPI_agent",uvm_component parent = null);
            super.new(name,parent);
        endfunction
        function void build_phase(uvm_phase phase);
            super.build_phase(phase);
            if(!uvm_config_db #(SPI_config_obj)::get(this,"","CFG",SPI_cfg))begin
                `uvm_fatal("bulid_phase","unable to get congiguration object")
            end
            sqr = SPI_sequencer::type_id::create("sqr",this);
            drv = SPI_driver::type_id::create("drv",this);
            mon = SPI_mon::type_id::create("mon",this);
            agt_ap = new("agt_ap",this);
        endfunction
        function void connect_phase(uvm_phase phase);
            super.connect_phase(phase);
            drv.SPI_vif = SPI_cfg.SPI_vif;
            mon.SPI_vif = SPI_cfg.SPI_vif;
            drv.seq_item_port.connect(sqr.seq_item_export);
            mon.mon_ap.connect(agt_ap);
        endfunction
    endclass
endpackage