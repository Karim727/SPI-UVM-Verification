module RAM (din,clk,rst_n,rx_valid,dout,tx_valid);

input      [9:0] din;
input            clk, rst_n, rx_valid;

output reg [7:0] dout;
output reg       tx_valid;

reg [7:0] MEM [255:0];

reg [7:0] Rd_Addr, Wr_Addr;

always @(posedge clk) begin
    if (~rst_n) begin
        dout <= 0;
        //tx_valid <= 0; <- BUG
        Rd_Addr <= 0;
        Wr_Addr <= 0;
    end
    else                                           
        if (rx_valid) begin
            case (din[9:8])
                2'b00 : Wr_Addr <= din[7:0]; // wr address
                2'b01 : MEM[Wr_Addr] <= din[7:0]; // wr data
                2'b10 : Rd_Addr <= din[7:0]; // rd address 
                2'b11 : dout <= MEM[Wr_Addr]; // rd data
                default : dout <= 0;
            endcase
        end
    tx_valid <= (din[9] && din[8] && rx_valid && rst_n)? 1'b1 : 1'b0;
end

endmodule