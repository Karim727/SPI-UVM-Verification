package RAM_shared_pkg;

endpackage