package RAM_shared_pkg;
    parameter RUNS = 1000;
endpackage