interface WRAPPER_if (clk);
  input clk;
  logic MOSI, SS_n, rst_n;
  logic MISO;
endinterface
