package WRAPPER_shared_pkg;
    paWRAPPEReter RUNS = 1000;
endpackage