package WRAPPER_shared_pkg;
    parameter RUNS = 1000;
    int count_ss_n = 0;
endpackage